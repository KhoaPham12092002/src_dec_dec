/* verilator lint_off UNUSED */
module single_cycle (
   input  logic           clk_i,
   input  logic           rst_ni,	
   input  logic  [W-1:0]  io_sw_i,

   output logic  [W-1:0]  pc_debug_o,
   output logic  [W-1:0]  io_lcd_o,
   output logic  [W-1:0]  io_ledg_o,
   output logic  [W-1:0]  io_ledr_o,
   output logic  [W-1:0]  io_hex0_o,
   output logic  [W-1:0]  io_hex1_o,
   output logic  [W-1:0]  io_hex2_o,
   output logic  [W-1:0]  io_hex3_o,
   output logic  [W-1:0]  io_hex4_o,
   output logic  [W-1:0]  io_hex5_o,
   output logic  [W-1:0]  io_hex6_o,
   output logic  [W-1:0]  io_hex7_o
);
parameter W = 32;
logic 	[W-1:0]  instr;
logic          	 br_eq;    
logic          	 br_lt; 
logic 	[2:0]    imm_gen_sel;  
logic 	[3:0]    alu_op;
logic          	 reg_wr_en;
logic          	 PC_sel;
logic          	 branch_u;
logic          	 dmem_wr;
logic          	 op_a_sel;
logic          	 op_b_sel;
logic 	[1:0]    wb_sel, fowardAE, fowardBE;
logic 	[W-1:0]  pc;
logic 	[W-1:0]  alu_data;
logic 	[W-1:0]  rs1_data, rs1_data_hazard;
logic 	[W-1:0]  rs2_data, rs2_data_hazard;
logic 	[W-1:0]  wb_data;
logic 	[W-1:0]  imm; 
logic 	[W-1:0]  operand_a;
logic 	[W-1:0]  operand_b;
logic 	[W-1:0]  ld_data;
logic 	[W-1:0]  digit9, digit8, digit7, digit6, digit5, digit4, digit3, digit2, digit1, digit0;
logic 	[3:0]    digit_sel;
logic 	[W-1:0]  digit_out;
logic   [W-1:0]  temp9, temp8, temp7, temp6, temp5, temp4, temp3, temp2, temp1, temp0;
logic            busy9, busy8, busy7, busy6, busy5, busy4, busy3, busy2, busy1, busy0;
logic            valid9, valid8, valid7, valid6, valid5, valid4, valid3, valid2, valid1, valid0;
logic            done9, done8, done7, done6, done5, done4, done3, done2, done1, done0;
logic		 start;
logic   [W-1:0]  pc_temp, instr_temp, pc_temp_temp, instr_temp_temp, rs1_data_temp, rs2_data_temp, imm_temp,
                 pc_temp_temp_temp, instr_temp_temp_temp, alu_data_temp, rs2_data_temp_temp,
                 pc_temp_temp_temp_temp, instr_temp_temp_temp_temp, alu_data_temp_temp, ld_data_temp,
		 instr_temp_temp_temp_temp_temp, wb_data_temp;
logic   [3:0]    alu_op_temp;
logic   [1:0]    wb_sel_temp, wb_sel_temp_temp, wb_sel_temp_temp_temp;
logic            reg_wr_en_temp, dmem_wr_temp, branch_u_temp, op_a_sel_temp, op_b_sel_temp, PC_sel_temp, reg_wr_en_temp_temp, dmem_wr_temp_temp, reg_wr_en_temp_temp_temp, hazard;
logic   [W-1:0] imm_hazard;
logic   [3:0]   alu_op_hazard;
logic   [1:0]   wb_sel_hazard;
logic           reg_wr_en_hazard, dmem_wr_hazard, branch_u_hazard, op_a_sel_hazard, op_b_sel_hazard, PC_sel_hazard;
logic           flushD;
logic           flushE;
logic           jump;
logic           PC_sel_br;
logic  [W-1:0]  PC_imm_addr;

assign flushD     = PC_sel_br;
assign flushE     = flushD|hazard;
assign pc_debug_o = pc;
assign PC_imm_addr = (instr_temp_temp[6:0] == 7'b1100111)? (imm_temp + operand_a):(imm_temp + pc_temp_temp);
assign PC_sel_br = jump & PC_sel_temp;

control_unit ctr_unit_block(
    .instr                        (instr_temp),
    .imm_gen_sel                  (imm_gen_sel),
    .alu_op                       (alu_op),
    .reg_wr_en                    (reg_wr_en),
    .PC_sel                       (PC_sel),
    .branch_u                     (branch_u),
    .dmem_wr                      (dmem_wr),
    .op_a_sel                     (op_a_sel),
    .op_b_sel                     (op_b_sel),
    .wb_sel                       (wb_sel)
);

hazard_unit hazard_unit_0 (
    .rs1_addr                     (instr_temp_temp[19:15]),
    .rs2_addr                     (instr_temp_temp[24:20]),
    .rdm_addr                     (instr_temp_temp_temp[11:7]),
    .rdw_addr                     (instr_temp_temp_temp_temp[11:7]),
    .rdt_addr                     (instr_temp_temp_temp_temp_temp[11:7]),
    .reg_wr_en_temp_temp          (reg_wr_en_temp_temp),
    .reg_wr_en_temp_temp_temp     (reg_wr_en_temp_temp_temp),
    .fowardAE                     (fowardAE),
    .fowardBE                     (fowardBE)
);

hazard_detect hazard_detect_0 (
   .IF_IDrs1_i                    (instr_temp[19:15]),
   .IF_IDrs2_i                    (instr_temp[24:20]),
   .ID_EXrd_i                     (instr_temp_temp[11:7]),
   .ID_EX_MemRead_i               (dmem_wr_temp),
   .hazard                        (hazard)
);

PC PC_block(
    .clk_i                        (clk_i),
    .rst_ni                       (rst_ni),
    .sel                          (PC_sel_br),
    .pc_imm                       (PC_imm_addr),
    .hazard                       (hazard),
    .pc_out                       (pc)
);

imem imem_block(
    .clk_i                        (clk_i),
    .rst_ni                       (rst_ni),
    .address                      (pc[13:0]),
    .data                         (instr)
);

reg_if_id reg_pipe_0(
    .clk_i                         (clk_i),
    .rst_ni                        (rst_ni),
    .flushD                        (flushD),
    .hazard                        (hazard),    
    .pc                            (pc),
    .instr                         (instr),
    .pc_temp                       (pc_temp),
    .instr_temp                    (instr_temp)
);

reg_32 regfile_block( 
    .clk_i                         (clk_i),
    .rst_ni                        (rst_ni),
    .addr_a                        (instr_temp[19:15]),
    .addr_b                        (instr_temp[24:20]),
    .addr_d                        (instr_temp_temp_temp_temp[11:7]),
    .data_d                        (wb_data),
    .wr_en_d                       (reg_wr_en_temp_temp_temp),
    .data_a                        (rs1_data),
    .data_b                        (rs2_data)
);

imm_gen immgen_block(
    .instr                         (instr_temp),      
    .imm_sel                       (imm_gen_sel),
    .imm                           (imm)
);

reg_id_ex reg_pipe_1(
    .clk_i                         (clk_i),
    .rst_ni                        (rst_ni),
    .flushE                        (flushE),
    .pc_temp                       (pc_temp),
    .instr_temp                    (instr_temp),
    .wb_sel                        (wb_sel),
    .reg_wr_en                     (reg_wr_en),
    .dmem_wr                       (dmem_wr),
    .rs1_data                      (rs1_data),
    .rs2_data                      (rs2_data),
    .alu_op                        (alu_op),
    .branch_u                      (branch_u),
    .op_a_sel                      (op_a_sel),
    .op_b_sel                      (op_b_sel),
    .imm                           (imm),
    .PC_sel                        (PC_sel),
    .pc_temp_temp                  (pc_temp_temp),
    .instr_temp_temp               (instr_temp_temp),
    .wb_sel_temp                   (wb_sel_temp),
    .reg_wr_en_temp                (reg_wr_en_temp),
    .dmem_wr_temp                  (dmem_wr_temp),
    .rs1_data_temp                 (rs1_data_temp),
    .rs2_data_temp                 (rs2_data_temp),
    .alu_op_temp                   (alu_op_temp),
    .branch_u_temp                 (branch_u_temp),
    .op_a_sel_temp                 (op_a_sel_temp),
    .op_b_sel_temp                 (op_b_sel_temp),
    .imm_temp                      (imm_temp),
    .PC_sel_temp                   (PC_sel_temp)
);	

branch_compare br_compare (
    .data_in_a                     (operand_a),
    .data_in_b                     (operand_b),
    .branch_unsigned               (branch_u_temp),
    .equal                         (br_eq),
    .lessthan                      (br_lt)
);

branch_control br_control (
    .instr                          (instr_temp_temp),
    .br_eq                          (br_eq),
    .br_lt                          (br_lt),
    .jump                           (jump)
);

mux_32bit_4x1 mux_hazard_0 (
    .a                              (rs1_data_temp),
    .b                              (wb_data),
    .c                              (alu_data_temp),
    .d                              (wb_data_temp),
    .sel                            (fowardAE),
    .out                            (rs1_data_hazard)
);

mux_32bit_4x1 mux_hazard_1 (
    .a                              (rs2_data_temp),
    .b                              (wb_data),
    .c                              (alu_data_temp),
    .d                              (wb_data_temp),
    .sel                            (fowardBE),
    .out                            (rs2_data_hazard)
);

mux_32bit mux_operand_a(
    .a                              (rs1_data_hazard),        
    .b                              (pc_temp_temp),
    .sel                            (op_a_sel_temp),
    .out                            (operand_a)
);

mux_32bit mux_operand_b(
    .a                              (rs2_data_hazard),        
    .b                              (imm_temp),
    .sel                            (op_b_sel_temp),
    .out                            (operand_b)
);

alu alu_block( 
    .in_alu_a                       (operand_a),
    .in_alu_b                       (operand_b),
    .alu_op                         (alu_op_temp),
    .branch_unsigned                (branch_u_temp),
    .out_alu                        (alu_data)
);

converter hex_to_dec (
    .clk                            (clk_i),
    .rst_n                          (rst_ni),
    .io_sw_i                        (io_sw_i),
    .result                         (rs1_data),
    .temp9                          (temp9),
    .temp8                          (temp8),
    .temp7                          (temp7),
    .temp6                          (temp6),
    .temp5                          (temp5),
    .temp4                          (temp4),
    .temp3                          (temp3),
    .temp2                          (temp2),
    .temp1                          (temp1),
    .temp0                          (temp0),
    .busy9                          (busy9),
    .busy8                          (busy8),
    .busy7                          (busy7),
    .busy6                          (busy6),
    .busy5                          (busy5),
    .busy4                          (busy4),
    .busy3                          (busy3),
    .busy2                          (busy2),
    .busy1                          (busy1),
    .busy0                          (busy0),
    .valid9                         (valid9),
    .valid8                         (valid8),
    .valid7                         (valid7),
    .valid6                         (valid6),
    .valid5                         (valid5),
    .valid4                         (valid4),
    .valid3                         (valid3),
    .valid2                         (valid2),
    .valid1                         (valid1),
    .valid0                         (valid0),
    .done9                          (done9),
    .done8                          (done8),
    .done7                          (done7),
    .done6                          (done6),
    .done5                          (done5),
    .done4                          (done4),
    .done3                          (done3),
    .done2                          (done2),
    .done1                          (done1),
    .done0                          (done0),
    .digit0                         (digit0),
    .digit1                         (digit1),
    .digit2                         (digit2),
    .digit3                         (digit3),
    .digit4                         (digit4),
    .digit5                         (digit5),
    .digit6                         (digit6),    
    .digit7                         (digit7),
    .digit8                         (digit8),
    .digit9                         (digit9)
);

reg_ex_mem reg_pipe_2(
    .clk_i                          (clk_i),
    .rst_ni                         (rst_ni),
    .pc_temp_temp                   (pc_temp_temp),
    .instr_temp_temp                (instr_temp_temp),
    .wb_sel_temp                    (wb_sel_temp),
    .reg_wr_en_temp                 (reg_wr_en_temp),
    .dmem_wr_temp                   (dmem_wr_temp),
    .alu_data                       (alu_data),
    .rs2_data_temp                  (rs2_data_hazard),
    .pc_temp_temp_temp              (pc_temp_temp_temp),
    .instr_temp_temp_temp           (instr_temp_temp_temp),
    .wb_sel_temp_temp               (wb_sel_temp_temp),
    .reg_wr_en_temp_temp            (reg_wr_en_temp_temp),
    .dmem_wr_temp_temp              (dmem_wr_temp_temp),
    .alu_data_temp                  (alu_data_temp),
    .rs2_data_temp_temp             (rs2_data_temp_temp)
);

dmem lsu_block(
    .clk_i                          (clk_i),        
    .rst_ni                         (rst_ni),
    .st_en                          (dmem_wr_temp_temp),
    .addr                           (alu_data_temp),    
    .unsigned_en_mem                (instr_temp_temp_temp[14]),
    .st_data                        (rs2_data_temp_temp),
    .sel_mod                        (instr_temp_temp_temp[13:12]),
    .io_sw_i                        (io_sw_i), 
    .ld_data                        (ld_data),    
    .io_lcd_o                       (io_lcd_o),    
    .io_ledg_o                      (io_ledg_o),    
    .io_ledr_o                      (io_ledr_o),    
    .io_hex0_o                      (io_hex0_o),
    .io_hex1_o                      (io_hex1_o),
    .io_hex2_o                      (io_hex2_o),
    .io_hex3_o                      (io_hex3_o),
    .io_hex4_o                      (io_hex4_o),
    .io_hex5_o                      (io_hex5_o),
    .io_hex6_o                      (io_hex6_o),
    .io_hex7_o                      (io_hex7_o)
);

mux_32bit_16x1 digit_sel_block(
    .a                              (digit0),
    .b                              (digit1),
    .c                              (digit2),
    .d                              (digit3),
    .e                              (digit4),
    .f                              (digit5),
    .g                              (digit6),
    .h                              (digit7),
    .j                              (digit8),
    .k                              (digit9),
    .l                              (32'b0),
    .m                              (32'b0),
    .n                              (32'b0),
    .q                              (32'b0),
    .r                              (32'b0),
    .s                              (32'b0),
    .sel                            (instr[31:28]),
    .out                            (digit_out)
);

reg_mem_wb reg_pipe_3(
    .clk_i                          (clk_i),
    .rst_ni                         (rst_ni),
    .pc_temp_temp_temp              (pc_temp_temp_temp),
    .instr_temp_temp_temp           (instr_temp_temp_temp),
    .wb_sel_temp_temp               (wb_sel_temp_temp),
    .alu_data_temp                  (alu_data_temp),
    .ld_data                        (ld_data),
    .reg_wr_en_temp_temp            (reg_wr_en_temp_temp),
    .pc_temp_temp_temp_temp         (pc_temp_temp_temp_temp),
    .instr_temp_temp_temp_temp      (instr_temp_temp_temp_temp),
    .wb_sel_temp_temp_temp          (wb_sel_temp_temp_temp),
    .alu_data_temp_temp             (alu_data_temp_temp),
    .ld_data_temp                   (ld_data_temp),
    .reg_wr_en_temp_temp_temp       (reg_wr_en_temp_temp_temp)
);

mux_32bit_4x1 wb_sel_block(
    .a                              (alu_data_temp_temp),
    .b                              (ld_data_temp),
    .c                              (pc_temp_temp_temp_temp),
    .d                              (digit_out),
    .sel                            (wb_sel_temp_temp_temp),
    .out                            (wb_data)
);

reg_rd reg_rd_0 (
    .clk_i                          (clk_i),
    .rst_ni                         (rst_ni),
    .instr_temp_temp_temp_temp      (instr_temp_temp_temp_temp),
    .wb_data                        (wb_data),
    .wb_data_temp                   (wb_data_temp),
    .instr_temp_temp_temp_temp_temp (instr_temp_temp_temp_temp_temp)
);

endmodule
